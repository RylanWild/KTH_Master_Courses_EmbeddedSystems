    Mac OS X            	   2   �      �                                      ATTR       �   �                      �      com.apple.quarantine q/0082;6578034b;prl_client_app; 