    Mac OS X            	   2   �      �                                      ATTR       �   �   0                  �     com.apple.lastuseddate#PS       �      com.apple.quarantine Q]xe    �Lg!    q/0082;6568f62e;prl_client_app; 