/*
@File    :   sigmoid_activation.sv
@Time    :   2023/11/24 10:05:57
@Author  :   Kevin Pettersson 
@Version :   1.0
@Contact :   kevinpet@kth.se
@License :   (C)Copyright 2023, Kevin Pettersson
@Desc    :   
*/


module sigmoid_activation (    
    input logic signed [7:0] input_data,
    
    output logic signed [7:0] output_data
);


always_comb begin
    case(input_data)
        8'b10000000 : output_data = 8'b00000000;
        8'b10000001 : output_data = 8'b00000000;
        8'b10000010 : output_data = 8'b00000000;
        8'b10000011 : output_data = 8'b00000000;
        8'b10000100 : output_data = 8'b00000000;
        8'b10000101 : output_data = 8'b00000000;
        8'b10000110 : output_data = 8'b00000000;
        8'b10000111 : output_data = 8'b00000000;
        8'b10001000 : output_data = 8'b00000000;
        8'b10001001 : output_data = 8'b00000000;
        8'b10001010 : output_data = 8'b00000000;
        8'b10001011 : output_data = 8'b00000000;
        8'b10001100 : output_data = 8'b00000000;
        8'b10001101 : output_data = 8'b00000000;
        8'b10001110 : output_data = 8'b00000000;
        8'b10001111 : output_data = 8'b00000000;
        8'b10010000 : output_data = 8'b00000000;
        8'b10010001 : output_data = 8'b00000000;
        8'b10010010 : output_data = 8'b00000000;
        8'b10010011 : output_data = 8'b00000001;
        8'b10010100 : output_data = 8'b00000001;
        8'b10010101 : output_data = 8'b00000001;
        8'b10010110 : output_data = 8'b00000001;
        8'b10010111 : output_data = 8'b00000001;
        8'b10011000 : output_data = 8'b00000001;
        8'b10011001 : output_data = 8'b00000001;
        8'b10011010 : output_data = 8'b00000001;
        8'b10011011 : output_data = 8'b00000001;
        8'b10011100 : output_data = 8'b00000001;
        8'b10011101 : output_data = 8'b00000001;
        8'b10011110 : output_data = 8'b00000001;
        8'b10011111 : output_data = 8'b00000001;
        8'b10100000 : output_data = 8'b00000001;
        8'b10100001 : output_data = 8'b00000001;
        8'b10100010 : output_data = 8'b00000001;
        8'b10100011 : output_data = 8'b00000001;
        8'b10100100 : output_data = 8'b00000001;
        8'b10100101 : output_data = 8'b00000001;
        8'b10100110 : output_data = 8'b00000001;
        8'b10100111 : output_data = 8'b00000001;
        8'b10101000 : output_data = 8'b00000001;
        8'b10101001 : output_data = 8'b00000001;
        8'b10101010 : output_data = 8'b00000010;
        8'b10101011 : output_data = 8'b00000010;
        8'b10101100 : output_data = 8'b00000010;
        8'b10101101 : output_data = 8'b00000010;
        8'b10101110 : output_data = 8'b00000010;
        8'b10101111 : output_data = 8'b00000010;
        8'b10110000 : output_data = 8'b00000010;
        8'b10110001 : output_data = 8'b00000010;
        8'b10110010 : output_data = 8'b00000010;
        8'b10110011 : output_data = 8'b00000010;
        8'b10110100 : output_data = 8'b00000010;
        8'b10110101 : output_data = 8'b00000010;
        8'b10110110 : output_data = 8'b00000010;
        8'b10110111 : output_data = 8'b00000010;
        8'b10111000 : output_data = 8'b00000011;
        8'b10111001 : output_data = 8'b00000011;
        8'b10111010 : output_data = 8'b00000011;
        8'b10111011 : output_data = 8'b00000011;
        8'b10111100 : output_data = 8'b00000011;
        8'b10111101 : output_data = 8'b00000011;
        8'b10111110 : output_data = 8'b00000011;
        8'b10111111 : output_data = 8'b00000011;
        8'b11000000 : output_data = 8'b00000011;
        8'b11000001 : output_data = 8'b00000011;
        8'b11000010 : output_data = 8'b00000100;
        8'b11000011 : output_data = 8'b00000100;
        8'b11000100 : output_data = 8'b00000100;
        8'b11000101 : output_data = 8'b00000100;
        8'b11000110 : output_data = 8'b00000100;
        8'b11000111 : output_data = 8'b00000100;
        8'b11001000 : output_data = 8'b00000100;
        8'b11001001 : output_data = 8'b00000100;
        8'b11001010 : output_data = 8'b00000100;
        8'b11001011 : output_data = 8'b00000101;
        8'b11001100 : output_data = 8'b00000101;
        8'b11001101 : output_data = 8'b00000101;
        8'b11001110 : output_data = 8'b00000101;
        8'b11001111 : output_data = 8'b00000101;
        8'b11010000 : output_data = 8'b00000101;
        8'b11010001 : output_data = 8'b00000101;
        8'b11010010 : output_data = 8'b00000110;
        8'b11010011 : output_data = 8'b00000110;
        8'b11010100 : output_data = 8'b00000110;
        8'b11010101 : output_data = 8'b00000110;
        8'b11010110 : output_data = 8'b00000110;
        8'b11010111 : output_data = 8'b00000110;
        8'b11011000 : output_data = 8'b00000111;
        8'b11011001 : output_data = 8'b00000111;
        8'b11011010 : output_data = 8'b00000111;
        8'b11011011 : output_data = 8'b00000111;
        8'b11011100 : output_data = 8'b00000111;
        8'b11011101 : output_data = 8'b00001000;
        8'b11011110 : output_data = 8'b00001000;
        8'b11011111 : output_data = 8'b00001000;
        8'b11100000 : output_data = 8'b00001000;
        8'b11100001 : output_data = 8'b00001000;
        8'b11100010 : output_data = 8'b00001001;
        8'b11100011 : output_data = 8'b00001001;
        8'b11100100 : output_data = 8'b00001001;
        8'b11100101 : output_data = 8'b00001001;
        8'b11100110 : output_data = 8'b00001001;
        8'b11100111 : output_data = 8'b00001010;
        8'b11101000 : output_data = 8'b00001010;
        8'b11101001 : output_data = 8'b00001010;
        8'b11101010 : output_data = 8'b00001010;
        8'b11101011 : output_data = 8'b00001010;
        8'b11101100 : output_data = 8'b00001011;
        8'b11101101 : output_data = 8'b00001011;
        8'b11101110 : output_data = 8'b00001011;
        8'b11101111 : output_data = 8'b00001011;
        8'b11110000 : output_data = 8'b00001100;
        8'b11110001 : output_data = 8'b00001100;
        8'b11110010 : output_data = 8'b00001100;
        8'b11110011 : output_data = 8'b00001100;
        8'b11110100 : output_data = 8'b00001101;
        8'b11110101 : output_data = 8'b00001101;
        8'b11110110 : output_data = 8'b00001101;
        8'b11110111 : output_data = 8'b00001101;
        8'b11111000 : output_data = 8'b00001110;
        8'b11111001 : output_data = 8'b00001110;
        8'b11111010 : output_data = 8'b00001110;
        8'b11111011 : output_data = 8'b00001110;
        8'b11111100 : output_data = 8'b00001111;
        8'b11111101 : output_data = 8'b00001111;
        8'b11111110 : output_data = 8'b00001111;
        8'b11111111 : output_data = 8'b00001111;
        8'b00000000 : output_data = 8'b00010000;
        8'b00000001 : output_data = 8'b00010000;
        8'b00000010 : output_data = 8'b00010000;
        8'b00000011 : output_data = 8'b00010000;
        8'b00000100 : output_data = 8'b00010000;
        8'b00000101 : output_data = 8'b00010001;
        8'b00000110 : output_data = 8'b00010001;
        8'b00000111 : output_data = 8'b00010001;
        8'b00001000 : output_data = 8'b00010001;
        8'b00001001 : output_data = 8'b00010010;
        8'b00001010 : output_data = 8'b00010010;
        8'b00001011 : output_data = 8'b00010010;
        8'b00001100 : output_data = 8'b00010010;
        8'b00001101 : output_data = 8'b00010011;
        8'b00001110 : output_data = 8'b00010011;
        8'b00001111 : output_data = 8'b00010011;
        8'b00010000 : output_data = 8'b00010011;
        8'b00010001 : output_data = 8'b00010100;
        8'b00010010 : output_data = 8'b00010100;
        8'b00010011 : output_data = 8'b00010100;
        8'b00010100 : output_data = 8'b00010100;
        8'b00010101 : output_data = 8'b00010101;
        8'b00010110 : output_data = 8'b00010101;
        8'b00010111 : output_data = 8'b00010101;
        8'b00011000 : output_data = 8'b00010101;
        8'b00011001 : output_data = 8'b00010101;
        8'b00011010 : output_data = 8'b00010110;
        8'b00011011 : output_data = 8'b00010110;
        8'b00011100 : output_data = 8'b00010110;
        8'b00011101 : output_data = 8'b00010110;
        8'b00011110 : output_data = 8'b00010110;
        8'b00011111 : output_data = 8'b00010111;
        8'b00100000 : output_data = 8'b00010111;
        8'b00100001 : output_data = 8'b00010111;
        8'b00100010 : output_data = 8'b00010111;
        8'b00100011 : output_data = 8'b00010111;
        8'b00100100 : output_data = 8'b00011000;
        8'b00100101 : output_data = 8'b00011000;
        8'b00100110 : output_data = 8'b00011000;
        8'b00100111 : output_data = 8'b00011000;
        8'b00101000 : output_data = 8'b00011000;
        8'b00101001 : output_data = 8'b00011001;
        8'b00101010 : output_data = 8'b00011001;
        8'b00101011 : output_data = 8'b00011001;
        8'b00101100 : output_data = 8'b00011001;
        8'b00101101 : output_data = 8'b00011001;
        8'b00101110 : output_data = 8'b00011001;
        8'b00101111 : output_data = 8'b00011010;
        8'b00110000 : output_data = 8'b00011010;
        8'b00110001 : output_data = 8'b00011010;
        8'b00110010 : output_data = 8'b00011010;
        8'b00110011 : output_data = 8'b00011010;
        8'b00110100 : output_data = 8'b00011010;
        8'b00110101 : output_data = 8'b00011010;
        8'b00110110 : output_data = 8'b00011011;
        8'b00110111 : output_data = 8'b00011011;
        8'b00111000 : output_data = 8'b00011011;
        8'b00111001 : output_data = 8'b00011011;
        8'b00111010 : output_data = 8'b00011011;
        8'b00111011 : output_data = 8'b00011011;
        8'b00111100 : output_data = 8'b00011011;
        8'b00111101 : output_data = 8'b00011011;
        8'b00111110 : output_data = 8'b00011011;
        8'b00111111 : output_data = 8'b00011100;
        8'b01000000 : output_data = 8'b00011100;
        8'b01000001 : output_data = 8'b00011100;
        8'b01000010 : output_data = 8'b00011100;
        8'b01000011 : output_data = 8'b00011100;
        8'b01000100 : output_data = 8'b00011100;
        8'b01000101 : output_data = 8'b00011100;
        8'b01000110 : output_data = 8'b00011100;
        8'b01000111 : output_data = 8'b00011100;
        8'b01001000 : output_data = 8'b00011100;
        8'b01001001 : output_data = 8'b00011101;
        8'b01001010 : output_data = 8'b00011101;
        8'b01001011 : output_data = 8'b00011101;
        8'b01001100 : output_data = 8'b00011101;
        8'b01001101 : output_data = 8'b00011101;
        8'b01001110 : output_data = 8'b00011101;
        8'b01001111 : output_data = 8'b00011101;
        8'b01010000 : output_data = 8'b00011101;
        8'b01010001 : output_data = 8'b00011101;
        8'b01010010 : output_data = 8'b00011101;
        8'b01010011 : output_data = 8'b00011101;
        8'b01010100 : output_data = 8'b00011101;
        8'b01010101 : output_data = 8'b00011101;
        8'b01010110 : output_data = 8'b00011101;
        8'b01010111 : output_data = 8'b00011110;
        8'b01011000 : output_data = 8'b00011110;
        8'b01011001 : output_data = 8'b00011110;
        8'b01011010 : output_data = 8'b00011110;
        8'b01011011 : output_data = 8'b00011110;
        8'b01011100 : output_data = 8'b00011110;
        8'b01011101 : output_data = 8'b00011110;
        8'b01011110 : output_data = 8'b00011110;
        8'b01011111 : output_data = 8'b00011110;
        8'b01100000 : output_data = 8'b00011110;
        8'b01100001 : output_data = 8'b00011110;
        8'b01100010 : output_data = 8'b00011110;
        8'b01100011 : output_data = 8'b00011110;
        8'b01100100 : output_data = 8'b00011110;
        8'b01100101 : output_data = 8'b00011110;
        8'b01100110 : output_data = 8'b00011110;
        8'b01100111 : output_data = 8'b00011110;
        8'b01101000 : output_data = 8'b00011110;
        8'b01101001 : output_data = 8'b00011110;
        8'b01101010 : output_data = 8'b00011110;
        8'b01101011 : output_data = 8'b00011110;
        8'b01101100 : output_data = 8'b00011110;
        8'b01101101 : output_data = 8'b00011110;
        8'b01101110 : output_data = 8'b00011111;
        8'b01101111 : output_data = 8'b00011111;
        8'b01110000 : output_data = 8'b00011111;
        8'b01110001 : output_data = 8'b00011111;
        8'b01110010 : output_data = 8'b00011111;
        8'b01110011 : output_data = 8'b00011111;
        8'b01110100 : output_data = 8'b00011111;
        8'b01110101 : output_data = 8'b00011111;
        8'b01110110 : output_data = 8'b00011111;
        8'b01110111 : output_data = 8'b00011111;
        8'b01111000 : output_data = 8'b00011111;
        8'b01111001 : output_data = 8'b00011111;
        8'b01111010 : output_data = 8'b00011111;
        8'b01111011 : output_data = 8'b00011111;
        8'b01111100 : output_data = 8'b00011111;
        8'b01111101 : output_data = 8'b00011111;
        8'b01111110 : output_data = 8'b00011111;
        8'b01111111 : output_data = 8'b00011111;
        default : output_data = 8'b00000000;
    endcase
end


endmodule