    Mac OS X            	   2   �      �                                      ATTR       �   �                      �      com.apple.quarantine q/0082;6568f62e;prl_client_app; 