    Mac OS X            	   2  #     U                                      ATTR      U  4  !                 4     com.apple.lastuseddate#PS      D   J  %com.apple.metadata:kMDItemWhereFroms   �  �  7com.apple.metadata:kMDLabel_tf3ulo4iwq7lwsunglwhmlkuem        >  com.apple.quarantine 4^xe    �>�1    bplist00�XHui Fengi i P h o n er�N N�                            '���#�g�g]��j�}hm�l�'��8�W����A��?H��q��ˎE������rvB����<��g��h��Ej�������z���7[e�c��N�K0��̝�����C�X�/����Ԣ��H��0�G�w���B]�iu��8v�)C8���ăT�{)X��ϧJ������i(.0�h2#�/s)�D����Q&��@B��n�%���o����� �CB��+�A�:~�"csQ~
��Ċ��6�#[D�y���F�W�3��*��'Z^>,Z[1�#knXS�yCn��~�a���=(�'˜̇��M�X��F�$jS��l �%���L���Qxn�_���0��-�̀�
'����*�������IE���U��O΂�W�у�q/0081;65785cfa;sharingd;D2094310-BAF2-4B94-A277-E5993172B419 