`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/09/25 05:54:26
// Design Name: 
// Module Name: weight
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package weight;
  
  parameter logic signed [7:0] weight_0 = 1;
  parameter logic signed [7:0] weight_1 = 2;
  parameter logic signed [7:0] weight_2 = 2;
  parameter logic signed [7:0] weight_3 = 2;
  parameter logic signed [7:0] weight_4 = 2;
  parameter logic signed [7:0] weight_5 = 1;
endpackage
