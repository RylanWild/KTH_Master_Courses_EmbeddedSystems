    Mac OS X            	   2  �                                           ATTR           �                       com.apple.lastuseddate#PS      0   H  com.apple.macl     x  i  7com.apple.metadata:kMDLabel_6r5l7e5tgj3mdhj6ygejexwizi     �      com.apple.quarantine �9xe    ��@/     �Z[�*H.��>Gl�� 5-ʾp�N��)q�f0��                                    ���V�������y��~���	���<���Fi�"��UD���B�5�n�}`��'������fY�J?�D�'��(�(I�C��!�"����� _��џO� �6��������&H!U��d�(��b���Kv���I��6rB�'=���*\�|0+i�x��Z���߬�$X;��@���0��u��F/�a�Vf���Պ���f�`lD�*(��V���n@�i�si��ݟ�^6�i��3�	��S��KB].��j�'��g�2�4�N�r(��@��0d0M �`?����3\�~5@�*���:�R��S�K�=�O�}γ�����tw7�$���25�5��6NK��*����{�kn�q/0082;6578079e;prl_client_app; 