    Mac OS X            	   2  �                                           ATTR                              J  %com.apple.metadata:kMDItemWhereFroms   V  �  7com.apple.metadata:kMDLabel_tf3ulo4iwq7lwsunglwhmlkuem     �   >  com.apple.quarantine bplist00�XHui Fengi i P h o n er�N N�                            '�b�!��d~�<�_���îu�Q [�N:�IN6�����NR԰�=�HL��Q�V�H���KQ ~�i���: }ʞ�.�M�1��qfyr�����7�E���Q�M.�T�Hu��,�����a��s/��f�K�̍I~wl�����9���J(�� ���B�l-�ց&-��␱K��n�c��v�Uł���~������@3��f|H�y ��D���z�����/�[��g[����û��c�|��+�R�و>k�|��Չ:���/���ǉ�`����ol)Kɛc���C��	�-���ƙ+�;Dj���8�ǵݵ��2��Y���z�uDDm�;�p��a�[��v�'�n�|>�c�ff��.�q/0081;65785d03;sharingd;BC833F23-3A4C-4E92-B807-6A122E44B136 