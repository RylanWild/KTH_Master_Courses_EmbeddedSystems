    Mac OS X            	   2  �                                           ATTR                              J  %com.apple.metadata:kMDItemWhereFroms   V  �  7com.apple.metadata:kMDLabel_tf3ulo4iwq7lwsunglwhmlkuem     �   >  com.apple.quarantine bplist00�XHui Fengi i P h o n er�N N�                            '��B�>�ٮ�B_C��g��Dt 쫐ȏw%�g Ro��ԛ,O��c.���yuG�������D��O��磨�`���4��f�[�@�E����rT��+~5r{F�����|]��J�J�3��.�`��h�4hr�1`A��?�λQ�L����Ǣ?��{�؊ٞD�E����A�8�qT�ؒ��3hǼ�/������^�mp#x��|��R�F�]�C��i��D�2�bSHR��P��WC V=��ꯘq6�3��%�p�>��ڰ���GQ��������:���q�U}�#��t�糵�x�P%�b6�8�?;�'m/�͉/��x$�R�R����Ux�!
Mȋ�?��|L/��%�v�i�I�ʆ���0�[m������
�"ͨUj�7q/0081;65785cef;sharingd;61F78C6A-A69C-4298-87B2-37F59568F454 